package pkg;
 
int number_of_transactions=20;
`include"trans.sv"
`include"gen.sv"
`include"drv.sv"
`include"wrmon.sv"
`include"rdmon.sv"
`include"rm.sv"
`include"sb.sv"
`include"env.sv"

endpackage
